library verilog;
use verilog.vl_types.all;
entity yusuf_gassaloglu_2020510034_HW1_a_vlg_sample_tst is
    port(
        clock           : in     vl_logic;
        count           : in     vl_logic;
        D0              : in     vl_logic;
        D1              : in     vl_logic;
        D2              : in     vl_logic;
        D3              : in     vl_logic;
        load            : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end yusuf_gassaloglu_2020510034_HW1_a_vlg_sample_tst;
