library verilog;
use verilog.vl_types.all;
entity yusuf_gassaloglu_2020510034_HW1_a is
    port(
        co              : out    vl_logic;
        count           : in     vl_logic;
        load            : in     vl_logic;
        D0              : in     vl_logic;
        clock           : in     vl_logic;
        D1              : in     vl_logic;
        D2              : in     vl_logic;
        D3              : in     vl_logic;
        Q0              : out    vl_logic;
        Q1              : out    vl_logic;
        Q2              : out    vl_logic;
        Q3              : out    vl_logic
    );
end yusuf_gassaloglu_2020510034_HW1_a;
