library verilog;
use verilog.vl_types.all;
entity yusuf_gassaloglu_2020510034_HW1_b_vlg_check_tst is
    port(
        carry           : in     vl_logic;
        q               : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end yusuf_gassaloglu_2020510034_HW1_b_vlg_check_tst;
