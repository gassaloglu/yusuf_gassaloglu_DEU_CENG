library verilog;
use verilog.vl_types.all;
entity \2020510034_Yusuf_group19_ALU\ is
    port(
        V               : out    vl_logic;
        Rs              : in     vl_logic_vector(3 downto 0);
        S2              : in     vl_logic_vector(3 downto 0);
        X               : in     vl_logic_vector(3 downto 0);
        Rd              : out    vl_logic_vector(3 downto 0)
    );
end \2020510034_Yusuf_group19_ALU\;
