library verilog;
use verilog.vl_types.all;
entity yusuf_gassaloglu_2020510034_HW1_a_vlg_check_tst is
    port(
        co              : in     vl_logic;
        Q0              : in     vl_logic;
        Q1              : in     vl_logic;
        Q2              : in     vl_logic;
        Q3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end yusuf_gassaloglu_2020510034_HW1_a_vlg_check_tst;
