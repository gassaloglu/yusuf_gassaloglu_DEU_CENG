library verilog;
use verilog.vl_types.all;
entity yusuf_gassaloglu_2020510034_HW1_a_vlg_vec_tst is
end yusuf_gassaloglu_2020510034_HW1_a_vlg_vec_tst;
