library verilog;
use verilog.vl_types.all;
entity yusuf_gassaloglu_2020510034_HW2_vlg_check_tst is
    port(
        ram_out         : in     vl_logic_vector(3 downto 0);
        rom_out         : in     vl_logic_vector(10 downto 0);
        sampler_rx      : in     vl_logic
    );
end yusuf_gassaloglu_2020510034_HW2_vlg_check_tst;
